//2022-7-19 反向器设计;


module inv(
	A,
	Y
	);
 	input A;
	output Y;

assign  Y=~A;

endmodule
